module BoomIOMSHR #(parameter id = 0)(
  input clock,
  input reset,

  Decouple.out io_req, //BoomDCacheReqST
  Decouple.in io_resp, //BoomDCacheRespST
  Decouple.in io_mem_access, //TLBundleA
  ValidSTIF.out io_mem_ack //TLBundleD
);
  
endmodule